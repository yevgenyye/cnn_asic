///////////////////////////////////////////////////////////////////////////////
// File Downloaded from http://www.nandland.com
///////////////////////////////////////////////////////////////////////////////
 `timescale 1 ns/10 ps 
//`include "carry_lookahead_adder.v"
 
module Huffman_enc_tb ();
 
  parameter W = 8;
  parameter C = 4;

  reg           clk     ;
  reg           rst     ;
  reg  [W-1:0]  d_in    ; // Huffman coded data
  reg  [C-1:0]  w_in    ;
  reg           en_in   ; // 
 
  wire [W-1:0]  d_out   ; // Encoded data
  wire          en_out  ; // 

  reg         init_end     ;

  integer     i,j;
 


localparam  B2_0   = 2'b00;    //W2_1 = 2;
localparam  B2_1   = 2'b01;    //W2_0 = 2;
localparam  B3_0   = 3'b100;   //W3_1 = 3;
localparam  B3_1   = 3'b101;   //W3_0 = 3;
localparam  B4_0   = 4'b1100;  //W4_1 = 4;
localparam  B4_1   = 4'b1101;  //W4_0 = 4;
localparam  B5_0   = 5'b11100; //W5_1 = 5;
localparam  B5_1   = 5'b11101; //W5_0 = 5;

localparam  B6_0   = 6'b111100;   //W6_1 = 6; 
localparam  B6_1   = 6'b111101;   //W6_0 = 6; 
localparam  B7_0   = 7'b1111100;  //W7_1 = 7; 
localparam  B7_1   = 7'b1111101;  //W7_0 = 7; 
localparam  B8_0   = 8'b11111100; //W8_1 = 8; 
localparam  B8_1   = 8'b11111101; //W8_0 = 8; 


  Huffman_enc  #(
    .W(W),
    .C(C)
    )
  DUT
  (
   .clk     (clk     ),
   .rst     (rst     ),
   .d_in    (d_in    ), // Huffman coded data
   .w_in    (w_in    ), 
   .en_in   (en_in   ), // 
   .d_out   (d_out   ), // Encoded data
   .en_out  (en_out  )  // 
   );

always 
begin
    clk = 1'b1; 
    #5; // high for 20 * timescale = 20 ns

    clk = 1'b0;
    #5; // low for 20 * timescale = 20 ns
end
 

   initial
     begin
           rst      <= 1'b1; 
           en_in    <= 0; 
       #10;
           rst   <= 1'b0; 
 
       #10;
       #10;
       #10;
 ////////////////////////////// operational part
        j= 0;
        #10;
        for (i = 0; i < 200; i = i + 1) 
          begin
            #10;
            j <= j + 1;
            en_in <= 1;
            $display("din(%h)= %h",i, d_in);
          end
         #10;
         en_in <= 0; 
 
         #100;
     end



 always @*
  case (j)
 
     1:  begin    d_in = { B2_0 , {(2){1'b0}} } ; w_in = 2; end // 1 byte 4x2
     2:  begin    d_in = { B2_1 , {(2){1'b0}} } ; w_in = 2; end //
     3:  begin    d_in = { B2_0 , {(2){1'b0}} } ; w_in = 2; end //
     4:  begin    d_in = { B2_1 , {(2){1'b0}} } ; w_in = 2; end //
     5:  begin    d_in = { B2_0 , {(2){1'b0}} } ; w_in = 2; end // 1 byte 4x2
     6:  begin    d_in = { B2_1 , {(2){1'b0}} } ; w_in = 2; end //
     7:  begin    d_in = { B2_0 , {(2){1'b0}} } ; w_in = 2; end //
     8:  begin    d_in = { B2_1 , {(2){1'b0}} } ; w_in = 2; end // 
     9:  begin    d_in = { B3_0 , {(3){1'b0}} } ; w_in = 3; end // 4 bytes 8x3
    10:  begin    d_in = { B3_1 , {(3){1'b0}} } ; w_in = 3; end //
    11:  begin    d_in = { B3_0 , {(3){1'b0}} } ; w_in = 3; end //
    12:  begin    d_in = { B3_1 , {(3){1'b0}} } ; w_in = 3; end //
    13:  begin    d_in = { B3_0 , {(3){1'b0}} } ; w_in = 3; end // 
    14:  begin    d_in = { B3_1 , {(3){1'b0}} } ; w_in = 3; end //
    15:  begin    d_in = { B3_0 , {(3){1'b0}} } ; w_in = 3; end //
    16:  begin    d_in = { B3_1 , {(3){1'b0}} } ; w_in = 3; end // 
 // 17:  begin    d_in = { }; //
 // 18:  begin    d_in = { }; //
 // 19:  begin    d_in = { }; //
 // 20:  begin    d_in = { }; //
 // 21:  begin    d_in = { }; //
 // 22:  begin    d_in = { }; //
 // 23:  begin    d_in = { }; // 
 // 24:  begin    d_in = { };
 // 25:  begin    d_in = { }; // 
 // 26:  begin    d_in = { }; //
 
  default:  d_in = 8'hFF;  
 endcase

endmodule // carry_lookahead_adder_tb